Library IEEE;
Use IEEE.Std_logic_1164.all;
Use IEEE.Std_logic_arith.all;
Use IEEE.Std_logic_unsigned.all;
entity divisor is
	Port( reloj: in std_logic;
			div_reloj : out std_logic);
end divisor;

architecture behavioral of divisor is
begin
	process (reloj)
		Constant N : integer := 16;
		variable cuenta : std_logic_vector (27 downto 0) := X"0000000";
		begin
			if rising_edge(reloj) then
				cuenta := cuenta + 1;
			end if;
			div_reloj <= cuenta(N);
	end process;
end behavioral;
--- Periodo de la señal de salida en función del valor N para un reloj = 50 MHZ
-- 27 – 5.37s, 26 – 2.68s, 25 – 1.34s, 24 – 671ms, 23 – 336ms
-- 22 – 168ms, 21 – 83.9ms, 20 – 41.9ms, 19 – 21ms, 18 – 10.5ms
-- 17 – 5.24ms, 16 – 2.62ms, 15 – 1.31ms, 14 – 655us, 13 – 320us
-- 12 – 164us, 11 – 81.9us, 10 – 41us, 9 – 20.5us, 8 – 10.2us
