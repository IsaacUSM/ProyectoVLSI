Library IEEE;
Use IEEE.Std_logic_1164.all;
Use IEEE.Std_logic_unsigned.all;
entity Teclado is
	Generic (FREQ_CLK: integer := 50_000_00);
	Port( CLK: IN STD_LOGIC;
			COLUMNAS: in std_logic_vector(3 downto 0);
			FILAS: out std_logic_vector(3 downto 0);
			reset: out std_logic;
			leftt:out std_logic;
			rightt:out std_logic;
			up:out std_logic;
			down:out std_logic;
			IND: out std_logic);
end Teclado;

architecture behavioral of Teclado is
	CONSTANT DELAY_1MS : INTEGER := (FREQ_CLK/1000)-1;
	CONSTANT DELAY_10MS : INTEGER := (FREQ_CLK/100)-1;
	SIGNAL CONTA_1MS: INTEGER RANGE 0 TO DELAY_1MS := 0;
	SIGNAL BANDERA: STD_LOGIC := '0';
	SIGNAL CONTA_10MS: INTEGER RANGE 0 TO DELAY_10MS := 0;
	SIGNAL BANDERA2 : STD_LOGIC := '0';
	SIGNAL BOT_D : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
	SIGNAL BOT_2 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
	SIGNAL BOT_4 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
	SIGNAL BOT_6 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
	SIGNAL BOT_8 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
	SIGNAL FILA_REG_S : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS=>'0');
	SIGNAL FILA : INTEGER RANGE 0 TO 3 := 0;
	SIGNAL IND_S : STD_LOGIC := '0';
	SIGNAL EDO : INTEGER RANGE 0 TO 1 := 0;
	BEGIN
		FILAS <= FILA_REG_S;
		--RETARDO 1 MS--
		PROCESS(CLK)
		BEGIN
			IF RISING_EDGE(CLK) THEN
				CONTA_1MS <= CONTA_1MS+1;
				BANDERA <= '0';
				IF CONTA_1MS = DELAY_1MS THEN
					CONTA_1MS <= 0;
					BANDERA <= '1';
				END IF;
			END IF;
		END PROCESS;
		----------------
		--RETARDO 10 MS--
		PROCESS(CLK)
		BEGIN
			IF RISING_EDGE(CLK) THEN
				CONTA_10MS <= CONTA_10MS+1;
				BANDERA2 <= '0';
				IF CONTA_10MS = DELAY_10MS THEN
					CONTA_10MS <= 0;
					BANDERA2 <= '1';
				END IF;
			END IF;
		END PROCESS;
		----------------
		--PROCESO EN LAS FILAS ----
		PROCESS(CLK, BANDERA2)
		BEGIN
			IF RISING_EDGE(CLK) AND BANDERA2 = '1' THEN
				FILA <= FILA+1;
				IF FILA = 3 THEN
					FILA <= 0;
				END IF;
			END IF;
		END PROCESS;
		WITH FILA SELECT
			FILA_REG_S <= 	"1000" WHEN 0,
								"0100" WHEN 1,
								"0010" WHEN 2,
								"0001" WHEN OTHERS;
		-------------------------------
		----------PROCESO EN EL TECLADO AL SELECCIONAR UN VALOR------------
		PROCESS(CLK,BANDERA)
		BEGIN
			IF RISING_EDGE(CLK) AND BANDERA = '1' THEN
				IF FILA_REG_S = "1000" THEN
					BOT_2 <= BOT_2(6 DOWNTO 0)&COLUMNAS(2);
				ELSIF FILA_REG_S = "0100" THEN
					BOT_4 <= BOT_4(6 DOWNTO 0)&COLUMNAS(3);
					BOT_6 <= BOT_6(6 DOWNTO 0)&COLUMNAS(1);
				ELSIF FILA_REG_S = "0010" THEN
					BOT_8 <= BOT_8(6 DOWNTO 0)&COLUMNAS(2);
				ELSIF FILA_REG_S = "0001" THEN
					BOT_D <= BOT_D(6 DOWNTO 0)&COLUMNAS(0);
				END IF;
			END IF;
		END PROCESS;
		----------------------------------------------------------------------------
		--SALIDA--
		PROCESS(CLK)
		BEGIN
			IF RISING_EDGE(CLK) THEN
				IF BOT_2 = "11111111" THEN 
					reset <= '0';
					leftt<= '0';
					rightt<= '0';
					up<= '1';
					down<= '0'; 
					IND_S <= '1';
				ELSIF BOT_4 = "11111111" THEN 
					reset <= '0';
					leftt<= '1';
					rightt<= '0';
					up<= '0';
					down<= '0'; 
					IND_S <= '1';
				ELSIF BOT_6 = "11111111" THEN 
					reset <= '0';
					leftt<= '0';
					rightt<= '1';
					up<= '0';
					down<= '0'; 
					IND_S <= '1';
				ELSIF BOT_8 = "11111111" THEN 
					reset <= '0';
					leftt<= '0';
					rightt<= '0';
					up<= '0';
					down<= '1'; 
					IND_S <= '1';
				ELSIF BOT_D = "11111111" THEN 
					reset <= '1';
					leftt<= '0';
					rightt<= '0';
					up<= '0';
					down<= '0'; 
					IND_S <= '1';
				ELSE 
					IND_S <= '0';
				END IF;
			END IF;
		END PROCESS;
		-----------------------------		
		--ACTIVACIÓN PARA LA BANDERA UN CICLO DE RELOJ--
		PROCESS(CLK)
		BEGIN
			IF RISING_EDGE(CLK) THEN
				IF EDO = 0 THEN
					IF IND_S = '1' THEN
						IND <= '1';
						EDO <= 1;
					ELSE
						EDO <= 0;
						IND <= '0';
					END IF;
				ELSE
					IF IND_S = '1' THEN
						EDO <= 1;
						IND <= '0';
					ELSE
						EDO <= 0;
					END IF;
				END IF;
			END IF;
		END PROCESS;
	--------------------------------------
END behavioral;